--
-- VHDL Architecture Display.vgaDataCreator.green
--
-- Created:
--          by - axel.amand.UNKNOWN (WE2330806)
--          at - 11:49:25 27.07.2022
--
-- using Mentor Graphics HDL Designer(TM) 2019.2 (Build 5)
--
ARCHITECTURE green OF vgaDataCreator IS
BEGIN
	pixelValue <= "010";
END ARCHITECTURE green;

