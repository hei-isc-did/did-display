--
-- VHDL Architecture Display_test.display_tb.test
--
-- Created:
--          by - zas.UNKNOWN (ZASE60F)
--          at - 13:44:09 11.07.2022
--
-- using Mentor Graphics HDL Designer(TM) 2019.4 (Build 4)
--
ARCHITECTURE test OF display_tb IS
BEGIN
END ARCHITECTURE test;

